LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux10to1 IS
	PORT ( S : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
			D : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			R0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R4 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R5 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R6 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R7 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			G : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			O : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END mux10to1;

--Mux que interliga a entrada DIN ou um registrador ao barramento BusWires!
ARCHITECTURE Behavior OF mux10to1 IS
	BEGIN
		PROCESS (S)
			BEGIN
				CASE S IS
					WHEN "1000000000" => O <= R0;
					WHEN "0100000000" => O <= R1;
					WHEN "0010000000" => O <= R2;
					WHEN "0001000000" => O <= R3;
					WHEN "0000100000" => O <= R4;
					WHEN "0000010000" => O <= R5;
					WHEN "0000001000" => O <= R6;
					WHEN "0000000100" => O <= R7;
					WHEN "0000000010" => O <= G;
					WHEN OTHERS => O <= D;
				END CASE;
		END PROCESS;
END Behavior;